// testeio.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module testeio (
		output wire [31:0] chrom_seg_0_export,              //              chrom_seg_0.export
		output wire [31:0] chrom_seg_1_export,              //              chrom_seg_1.export
		output wire [31:0] chrom_seg_10_export,             //             chrom_seg_10.export
		output wire [31:0] chrom_seg_11_export,             //             chrom_seg_11.export
		output wire [31:0] chrom_seg_12_export,             //             chrom_seg_12.export
		output wire [31:0] chrom_seg_13_export,             //             chrom_seg_13.export
		output wire [31:0] chrom_seg_14_export,             //             chrom_seg_14.export
		output wire [31:0] chrom_seg_15_export,             //             chrom_seg_15.export
		output wire [31:0] chrom_seg_16_export,             //             chrom_seg_16.export
		output wire [31:0] chrom_seg_17_export,             //             chrom_seg_17.export
		output wire [31:0] chrom_seg_18_export,             //             chrom_seg_18.export
		output wire [31:0] chrom_seg_19_export,             //             chrom_seg_19.export
		output wire [31:0] chrom_seg_2_export,              //              chrom_seg_2.export
		output wire [31:0] chrom_seg_20_export,             //             chrom_seg_20.export
		output wire [31:0] chrom_seg_21_export,             //             chrom_seg_21.export
		output wire [31:0] chrom_seg_22_export,             //             chrom_seg_22.export
		output wire [31:0] chrom_seg_23_export,             //             chrom_seg_23.export
		output wire [31:0] chrom_seg_24_export,             //             chrom_seg_24.export
		output wire [31:0] chrom_seg_25_export,             //             chrom_seg_25.export
		output wire [31:0] chrom_seg_26_export,             //             chrom_seg_26.export
		output wire [31:0] chrom_seg_27_export,             //             chrom_seg_27.export
		output wire [31:0] chrom_seg_28_export,             //             chrom_seg_28.export
		output wire [31:0] chrom_seg_29_export,             //             chrom_seg_29.export
		output wire [31:0] chrom_seg_3_export,              //              chrom_seg_3.export
		output wire [31:0] chrom_seg_30_export,             //             chrom_seg_30.export
		output wire [31:0] chrom_seg_4_export,              //              chrom_seg_4.export
		output wire [31:0] chrom_seg_5_export,              //              chrom_seg_5.export
		output wire [31:0] chrom_seg_6_export,              //              chrom_seg_6.export
		output wire [31:0] chrom_seg_7_export,              //              chrom_seg_7.export
		output wire [31:0] chrom_seg_8_export,              //              chrom_seg_8.export
		output wire [31:0] chrom_seg_9_export,              //              chrom_seg_9.export
		input  wire        clk_clk,                         //                      clk.clk
		input  wire [14:0] correct_mem_s2_address,          //           correct_mem_s2.address
		input  wire        correct_mem_s2_chipselect,       //                         .chipselect
		input  wire        correct_mem_s2_clken,            //                         .clken
		input  wire        correct_mem_s2_write,            //                         .write
		output wire [31:0] correct_mem_s2_readdata,         //                         .readdata
		input  wire [31:0] correct_mem_s2_writedata,        //                         .writedata
		input  wire [3:0]  correct_mem_s2_byteenable,       //                         .byteenable
		input  wire        done_processing_chrom_export,    //    done_processing_chrom.export
		output wire        done_processing_feedback_export, // done_processing_feedback.export
		input  wire [31:0] error_sum_0_export,              //              error_sum_0.export
		input  wire [31:0] error_sum_1_export,              //              error_sum_1.export
		input  wire [31:0] error_sum_2_export,              //              error_sum_2.export
		input  wire [31:0] error_sum_3_export,              //              error_sum_3.export
		input  wire [31:0] error_sum_4_export,              //              error_sum_4.export
		input  wire [31:0] error_sum_5_export,              //              error_sum_5.export
		input  wire [31:0] error_sum_6_export,              //              error_sum_6.export
		input  wire [31:0] error_sum_7_export,              //              error_sum_7.export
		output wire [31:0] expected_output_0_export,        //        expected_output_0.export
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //                   hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //                         .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //                         .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //                         .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //                         .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //                         .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //                         .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //                         .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //                         .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //                         .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //                         .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //                         .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //                         .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //                         .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //                         .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //                         .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //                         .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //                         .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //                         .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //                         .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //                         .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //                         .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //                         .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //                         .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //                         .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //                         .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //                         .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //                         .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //                         .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //                         .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //                         .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //                         .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,     //                         .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //                         .hps_io_uart0_inst_TX
		output wire [31:0] input_sequence_0_export,         //         input_sequence_0.export
		input  wire [14:0] mem_s2_address,                  //                   mem_s2.address
		input  wire        mem_s2_chipselect,               //                         .chipselect
		input  wire        mem_s2_clken,                    //                         .clken
		input  wire        mem_s2_write,                    //                         .write
		output wire [31:0] mem_s2_readdata,                 //                         .readdata
		input  wire [31:0] mem_s2_writedata,                //                         .writedata
		input  wire [3:0]  mem_s2_byteenable,               //                         .byteenable
		output wire [14:0] memory_mem_a,                    //                   memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                         .mem_ba
		output wire        memory_mem_ck,                   //                         .mem_ck
		output wire        memory_mem_ck_n,                 //                         .mem_ck_n
		output wire        memory_mem_cke,                  //                         .mem_cke
		output wire        memory_mem_cs_n,                 //                         .mem_cs_n
		output wire        memory_mem_ras_n,                //                         .mem_ras_n
		output wire        memory_mem_cas_n,                //                         .mem_cas_n
		output wire        memory_mem_we_n,                 //                         .mem_we_n
		output wire        memory_mem_reset_n,              //                         .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //                         .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //                         .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //                         .mem_dqs_n
		output wire        memory_mem_odt,                  //                         .mem_odt
		output wire [3:0]  memory_mem_dm,                   //                         .mem_dm
		input  wire        memory_oct_rzqin,                //                         .oct_rzqin
		input  wire [31:0] nextsample_export,               //               nextsample.export
		output wire [31:0] preparingnextsample_export,      //      preparingnextsample.export
		input  wire        ready_to_process_export,         //         ready_to_process.export
		input  wire        reset_reset_n,                   //                    reset.reset_n
		output wire [31:0] sampleindex_export,              //              sampleindex.export
		output wire [31:0] sequences_to_process_export,     //     sequences_to_process.export
		output wire        start_processing_chrom_export,   //   start_processing_chrom.export
		output wire [31:0] valid_output_0_export,           //           valid_output_0.export
		output wire [31:0] writesample_export               //              writesample.export
	);

	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                          // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                            // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                            // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                              // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                           // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                            // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                              // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                          // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                           // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                           // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                           // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                           // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                            // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                          // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                          // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                             // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                           // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                           // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                           // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                          // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                           // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                           // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                            // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                             // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                              // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                           // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                          // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire         mm_interconnect_0_chrom_seg_0_s1_chipselect;              // mm_interconnect_0:chrom_seg_0_s1_chipselect -> chrom_seg_0:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_0_s1_readdata;                // chrom_seg_0:readdata -> mm_interconnect_0:chrom_seg_0_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_0_s1_address;                 // mm_interconnect_0:chrom_seg_0_s1_address -> chrom_seg_0:address
	wire         mm_interconnect_0_chrom_seg_0_s1_write;                   // mm_interconnect_0:chrom_seg_0_s1_write -> chrom_seg_0:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_0_s1_writedata;               // mm_interconnect_0:chrom_seg_0_s1_writedata -> chrom_seg_0:writedata
	wire         mm_interconnect_0_chrom_seg_1_s1_chipselect;              // mm_interconnect_0:chrom_seg_1_s1_chipselect -> chrom_seg_1:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_1_s1_readdata;                // chrom_seg_1:readdata -> mm_interconnect_0:chrom_seg_1_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_1_s1_address;                 // mm_interconnect_0:chrom_seg_1_s1_address -> chrom_seg_1:address
	wire         mm_interconnect_0_chrom_seg_1_s1_write;                   // mm_interconnect_0:chrom_seg_1_s1_write -> chrom_seg_1:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_1_s1_writedata;               // mm_interconnect_0:chrom_seg_1_s1_writedata -> chrom_seg_1:writedata
	wire         mm_interconnect_0_chrom_seg_2_s1_chipselect;              // mm_interconnect_0:chrom_seg_2_s1_chipselect -> chrom_seg_2:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_2_s1_readdata;                // chrom_seg_2:readdata -> mm_interconnect_0:chrom_seg_2_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_2_s1_address;                 // mm_interconnect_0:chrom_seg_2_s1_address -> chrom_seg_2:address
	wire         mm_interconnect_0_chrom_seg_2_s1_write;                   // mm_interconnect_0:chrom_seg_2_s1_write -> chrom_seg_2:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_2_s1_writedata;               // mm_interconnect_0:chrom_seg_2_s1_writedata -> chrom_seg_2:writedata
	wire         mm_interconnect_0_chrom_seg_3_s1_chipselect;              // mm_interconnect_0:chrom_seg_3_s1_chipselect -> chrom_seg_3:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_3_s1_readdata;                // chrom_seg_3:readdata -> mm_interconnect_0:chrom_seg_3_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_3_s1_address;                 // mm_interconnect_0:chrom_seg_3_s1_address -> chrom_seg_3:address
	wire         mm_interconnect_0_chrom_seg_3_s1_write;                   // mm_interconnect_0:chrom_seg_3_s1_write -> chrom_seg_3:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_3_s1_writedata;               // mm_interconnect_0:chrom_seg_3_s1_writedata -> chrom_seg_3:writedata
	wire         mm_interconnect_0_chrom_seg_4_s1_chipselect;              // mm_interconnect_0:chrom_seg_4_s1_chipselect -> chrom_seg_4:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_4_s1_readdata;                // chrom_seg_4:readdata -> mm_interconnect_0:chrom_seg_4_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_4_s1_address;                 // mm_interconnect_0:chrom_seg_4_s1_address -> chrom_seg_4:address
	wire         mm_interconnect_0_chrom_seg_4_s1_write;                   // mm_interconnect_0:chrom_seg_4_s1_write -> chrom_seg_4:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_4_s1_writedata;               // mm_interconnect_0:chrom_seg_4_s1_writedata -> chrom_seg_4:writedata
	wire         mm_interconnect_0_chrom_seg_5_s1_chipselect;              // mm_interconnect_0:chrom_seg_5_s1_chipselect -> chrom_seg_5:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_5_s1_readdata;                // chrom_seg_5:readdata -> mm_interconnect_0:chrom_seg_5_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_5_s1_address;                 // mm_interconnect_0:chrom_seg_5_s1_address -> chrom_seg_5:address
	wire         mm_interconnect_0_chrom_seg_5_s1_write;                   // mm_interconnect_0:chrom_seg_5_s1_write -> chrom_seg_5:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_5_s1_writedata;               // mm_interconnect_0:chrom_seg_5_s1_writedata -> chrom_seg_5:writedata
	wire         mm_interconnect_0_chrom_seg_6_s1_chipselect;              // mm_interconnect_0:chrom_seg_6_s1_chipselect -> chrom_seg_6:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_6_s1_readdata;                // chrom_seg_6:readdata -> mm_interconnect_0:chrom_seg_6_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_6_s1_address;                 // mm_interconnect_0:chrom_seg_6_s1_address -> chrom_seg_6:address
	wire         mm_interconnect_0_chrom_seg_6_s1_write;                   // mm_interconnect_0:chrom_seg_6_s1_write -> chrom_seg_6:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_6_s1_writedata;               // mm_interconnect_0:chrom_seg_6_s1_writedata -> chrom_seg_6:writedata
	wire         mm_interconnect_0_chrom_seg_7_s1_chipselect;              // mm_interconnect_0:chrom_seg_7_s1_chipselect -> chrom_seg_7:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_7_s1_readdata;                // chrom_seg_7:readdata -> mm_interconnect_0:chrom_seg_7_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_7_s1_address;                 // mm_interconnect_0:chrom_seg_7_s1_address -> chrom_seg_7:address
	wire         mm_interconnect_0_chrom_seg_7_s1_write;                   // mm_interconnect_0:chrom_seg_7_s1_write -> chrom_seg_7:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_7_s1_writedata;               // mm_interconnect_0:chrom_seg_7_s1_writedata -> chrom_seg_7:writedata
	wire         mm_interconnect_0_chrom_seg_8_s1_chipselect;              // mm_interconnect_0:chrom_seg_8_s1_chipselect -> chrom_seg_8:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_8_s1_readdata;                // chrom_seg_8:readdata -> mm_interconnect_0:chrom_seg_8_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_8_s1_address;                 // mm_interconnect_0:chrom_seg_8_s1_address -> chrom_seg_8:address
	wire         mm_interconnect_0_chrom_seg_8_s1_write;                   // mm_interconnect_0:chrom_seg_8_s1_write -> chrom_seg_8:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_8_s1_writedata;               // mm_interconnect_0:chrom_seg_8_s1_writedata -> chrom_seg_8:writedata
	wire         mm_interconnect_0_chrom_seg_9_s1_chipselect;              // mm_interconnect_0:chrom_seg_9_s1_chipselect -> chrom_seg_9:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_9_s1_readdata;                // chrom_seg_9:readdata -> mm_interconnect_0:chrom_seg_9_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_9_s1_address;                 // mm_interconnect_0:chrom_seg_9_s1_address -> chrom_seg_9:address
	wire         mm_interconnect_0_chrom_seg_9_s1_write;                   // mm_interconnect_0:chrom_seg_9_s1_write -> chrom_seg_9:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_9_s1_writedata;               // mm_interconnect_0:chrom_seg_9_s1_writedata -> chrom_seg_9:writedata
	wire         mm_interconnect_0_chrom_seg_10_s1_chipselect;             // mm_interconnect_0:chrom_seg_10_s1_chipselect -> chrom_seg_10:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_10_s1_readdata;               // chrom_seg_10:readdata -> mm_interconnect_0:chrom_seg_10_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_10_s1_address;                // mm_interconnect_0:chrom_seg_10_s1_address -> chrom_seg_10:address
	wire         mm_interconnect_0_chrom_seg_10_s1_write;                  // mm_interconnect_0:chrom_seg_10_s1_write -> chrom_seg_10:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_10_s1_writedata;              // mm_interconnect_0:chrom_seg_10_s1_writedata -> chrom_seg_10:writedata
	wire         mm_interconnect_0_chrom_seg_11_s1_chipselect;             // mm_interconnect_0:chrom_seg_11_s1_chipselect -> chrom_seg_11:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_11_s1_readdata;               // chrom_seg_11:readdata -> mm_interconnect_0:chrom_seg_11_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_11_s1_address;                // mm_interconnect_0:chrom_seg_11_s1_address -> chrom_seg_11:address
	wire         mm_interconnect_0_chrom_seg_11_s1_write;                  // mm_interconnect_0:chrom_seg_11_s1_write -> chrom_seg_11:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_11_s1_writedata;              // mm_interconnect_0:chrom_seg_11_s1_writedata -> chrom_seg_11:writedata
	wire         mm_interconnect_0_chrom_seg_12_s1_chipselect;             // mm_interconnect_0:chrom_seg_12_s1_chipselect -> chrom_seg_12:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_12_s1_readdata;               // chrom_seg_12:readdata -> mm_interconnect_0:chrom_seg_12_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_12_s1_address;                // mm_interconnect_0:chrom_seg_12_s1_address -> chrom_seg_12:address
	wire         mm_interconnect_0_chrom_seg_12_s1_write;                  // mm_interconnect_0:chrom_seg_12_s1_write -> chrom_seg_12:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_12_s1_writedata;              // mm_interconnect_0:chrom_seg_12_s1_writedata -> chrom_seg_12:writedata
	wire         mm_interconnect_0_chrom_seg_13_s1_chipselect;             // mm_interconnect_0:chrom_seg_13_s1_chipselect -> chrom_seg_13:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_13_s1_readdata;               // chrom_seg_13:readdata -> mm_interconnect_0:chrom_seg_13_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_13_s1_address;                // mm_interconnect_0:chrom_seg_13_s1_address -> chrom_seg_13:address
	wire         mm_interconnect_0_chrom_seg_13_s1_write;                  // mm_interconnect_0:chrom_seg_13_s1_write -> chrom_seg_13:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_13_s1_writedata;              // mm_interconnect_0:chrom_seg_13_s1_writedata -> chrom_seg_13:writedata
	wire         mm_interconnect_0_chrom_seg_14_s1_chipselect;             // mm_interconnect_0:chrom_seg_14_s1_chipselect -> chrom_seg_14:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_14_s1_readdata;               // chrom_seg_14:readdata -> mm_interconnect_0:chrom_seg_14_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_14_s1_address;                // mm_interconnect_0:chrom_seg_14_s1_address -> chrom_seg_14:address
	wire         mm_interconnect_0_chrom_seg_14_s1_write;                  // mm_interconnect_0:chrom_seg_14_s1_write -> chrom_seg_14:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_14_s1_writedata;              // mm_interconnect_0:chrom_seg_14_s1_writedata -> chrom_seg_14:writedata
	wire         mm_interconnect_0_chrom_seg_15_s1_chipselect;             // mm_interconnect_0:chrom_seg_15_s1_chipselect -> chrom_seg_15:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_15_s1_readdata;               // chrom_seg_15:readdata -> mm_interconnect_0:chrom_seg_15_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_15_s1_address;                // mm_interconnect_0:chrom_seg_15_s1_address -> chrom_seg_15:address
	wire         mm_interconnect_0_chrom_seg_15_s1_write;                  // mm_interconnect_0:chrom_seg_15_s1_write -> chrom_seg_15:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_15_s1_writedata;              // mm_interconnect_0:chrom_seg_15_s1_writedata -> chrom_seg_15:writedata
	wire         mm_interconnect_0_chrom_seg_16_s1_chipselect;             // mm_interconnect_0:chrom_seg_16_s1_chipselect -> chrom_seg_16:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_16_s1_readdata;               // chrom_seg_16:readdata -> mm_interconnect_0:chrom_seg_16_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_16_s1_address;                // mm_interconnect_0:chrom_seg_16_s1_address -> chrom_seg_16:address
	wire         mm_interconnect_0_chrom_seg_16_s1_write;                  // mm_interconnect_0:chrom_seg_16_s1_write -> chrom_seg_16:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_16_s1_writedata;              // mm_interconnect_0:chrom_seg_16_s1_writedata -> chrom_seg_16:writedata
	wire         mm_interconnect_0_chrom_seg_17_s1_chipselect;             // mm_interconnect_0:chrom_seg_17_s1_chipselect -> chrom_seg_17:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_17_s1_readdata;               // chrom_seg_17:readdata -> mm_interconnect_0:chrom_seg_17_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_17_s1_address;                // mm_interconnect_0:chrom_seg_17_s1_address -> chrom_seg_17:address
	wire         mm_interconnect_0_chrom_seg_17_s1_write;                  // mm_interconnect_0:chrom_seg_17_s1_write -> chrom_seg_17:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_17_s1_writedata;              // mm_interconnect_0:chrom_seg_17_s1_writedata -> chrom_seg_17:writedata
	wire         mm_interconnect_0_chrom_seg_18_s1_chipselect;             // mm_interconnect_0:chrom_seg_18_s1_chipselect -> chrom_seg_18:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_18_s1_readdata;               // chrom_seg_18:readdata -> mm_interconnect_0:chrom_seg_18_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_18_s1_address;                // mm_interconnect_0:chrom_seg_18_s1_address -> chrom_seg_18:address
	wire         mm_interconnect_0_chrom_seg_18_s1_write;                  // mm_interconnect_0:chrom_seg_18_s1_write -> chrom_seg_18:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_18_s1_writedata;              // mm_interconnect_0:chrom_seg_18_s1_writedata -> chrom_seg_18:writedata
	wire         mm_interconnect_0_chrom_seg_19_s1_chipselect;             // mm_interconnect_0:chrom_seg_19_s1_chipselect -> chrom_seg_19:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_19_s1_readdata;               // chrom_seg_19:readdata -> mm_interconnect_0:chrom_seg_19_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_19_s1_address;                // mm_interconnect_0:chrom_seg_19_s1_address -> chrom_seg_19:address
	wire         mm_interconnect_0_chrom_seg_19_s1_write;                  // mm_interconnect_0:chrom_seg_19_s1_write -> chrom_seg_19:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_19_s1_writedata;              // mm_interconnect_0:chrom_seg_19_s1_writedata -> chrom_seg_19:writedata
	wire         mm_interconnect_0_chrom_seg_20_s1_chipselect;             // mm_interconnect_0:chrom_seg_20_s1_chipselect -> chrom_seg_20:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_20_s1_readdata;               // chrom_seg_20:readdata -> mm_interconnect_0:chrom_seg_20_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_20_s1_address;                // mm_interconnect_0:chrom_seg_20_s1_address -> chrom_seg_20:address
	wire         mm_interconnect_0_chrom_seg_20_s1_write;                  // mm_interconnect_0:chrom_seg_20_s1_write -> chrom_seg_20:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_20_s1_writedata;              // mm_interconnect_0:chrom_seg_20_s1_writedata -> chrom_seg_20:writedata
	wire         mm_interconnect_0_chrom_seg_21_s1_chipselect;             // mm_interconnect_0:chrom_seg_21_s1_chipselect -> chrom_seg_21:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_21_s1_readdata;               // chrom_seg_21:readdata -> mm_interconnect_0:chrom_seg_21_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_21_s1_address;                // mm_interconnect_0:chrom_seg_21_s1_address -> chrom_seg_21:address
	wire         mm_interconnect_0_chrom_seg_21_s1_write;                  // mm_interconnect_0:chrom_seg_21_s1_write -> chrom_seg_21:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_21_s1_writedata;              // mm_interconnect_0:chrom_seg_21_s1_writedata -> chrom_seg_21:writedata
	wire         mm_interconnect_0_chrom_seg_22_s1_chipselect;             // mm_interconnect_0:chrom_seg_22_s1_chipselect -> chrom_seg_22:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_22_s1_readdata;               // chrom_seg_22:readdata -> mm_interconnect_0:chrom_seg_22_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_22_s1_address;                // mm_interconnect_0:chrom_seg_22_s1_address -> chrom_seg_22:address
	wire         mm_interconnect_0_chrom_seg_22_s1_write;                  // mm_interconnect_0:chrom_seg_22_s1_write -> chrom_seg_22:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_22_s1_writedata;              // mm_interconnect_0:chrom_seg_22_s1_writedata -> chrom_seg_22:writedata
	wire         mm_interconnect_0_chrom_seg_23_s1_chipselect;             // mm_interconnect_0:chrom_seg_23_s1_chipselect -> chrom_seg_23:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_23_s1_readdata;               // chrom_seg_23:readdata -> mm_interconnect_0:chrom_seg_23_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_23_s1_address;                // mm_interconnect_0:chrom_seg_23_s1_address -> chrom_seg_23:address
	wire         mm_interconnect_0_chrom_seg_23_s1_write;                  // mm_interconnect_0:chrom_seg_23_s1_write -> chrom_seg_23:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_23_s1_writedata;              // mm_interconnect_0:chrom_seg_23_s1_writedata -> chrom_seg_23:writedata
	wire         mm_interconnect_0_chrom_seg_24_s1_chipselect;             // mm_interconnect_0:chrom_seg_24_s1_chipselect -> chrom_seg_24:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_24_s1_readdata;               // chrom_seg_24:readdata -> mm_interconnect_0:chrom_seg_24_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_24_s1_address;                // mm_interconnect_0:chrom_seg_24_s1_address -> chrom_seg_24:address
	wire         mm_interconnect_0_chrom_seg_24_s1_write;                  // mm_interconnect_0:chrom_seg_24_s1_write -> chrom_seg_24:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_24_s1_writedata;              // mm_interconnect_0:chrom_seg_24_s1_writedata -> chrom_seg_24:writedata
	wire         mm_interconnect_0_chrom_seg_25_s1_chipselect;             // mm_interconnect_0:chrom_seg_25_s1_chipselect -> chrom_seg_25:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_25_s1_readdata;               // chrom_seg_25:readdata -> mm_interconnect_0:chrom_seg_25_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_25_s1_address;                // mm_interconnect_0:chrom_seg_25_s1_address -> chrom_seg_25:address
	wire         mm_interconnect_0_chrom_seg_25_s1_write;                  // mm_interconnect_0:chrom_seg_25_s1_write -> chrom_seg_25:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_25_s1_writedata;              // mm_interconnect_0:chrom_seg_25_s1_writedata -> chrom_seg_25:writedata
	wire         mm_interconnect_0_chrom_seg_26_s1_chipselect;             // mm_interconnect_0:chrom_seg_26_s1_chipselect -> chrom_seg_26:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_26_s1_readdata;               // chrom_seg_26:readdata -> mm_interconnect_0:chrom_seg_26_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_26_s1_address;                // mm_interconnect_0:chrom_seg_26_s1_address -> chrom_seg_26:address
	wire         mm_interconnect_0_chrom_seg_26_s1_write;                  // mm_interconnect_0:chrom_seg_26_s1_write -> chrom_seg_26:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_26_s1_writedata;              // mm_interconnect_0:chrom_seg_26_s1_writedata -> chrom_seg_26:writedata
	wire         mm_interconnect_0_chrom_seg_27_s1_chipselect;             // mm_interconnect_0:chrom_seg_27_s1_chipselect -> chrom_seg_27:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_27_s1_readdata;               // chrom_seg_27:readdata -> mm_interconnect_0:chrom_seg_27_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_27_s1_address;                // mm_interconnect_0:chrom_seg_27_s1_address -> chrom_seg_27:address
	wire         mm_interconnect_0_chrom_seg_27_s1_write;                  // mm_interconnect_0:chrom_seg_27_s1_write -> chrom_seg_27:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_27_s1_writedata;              // mm_interconnect_0:chrom_seg_27_s1_writedata -> chrom_seg_27:writedata
	wire         mm_interconnect_0_chrom_seg_28_s1_chipselect;             // mm_interconnect_0:chrom_seg_28_s1_chipselect -> chrom_seg_28:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_28_s1_readdata;               // chrom_seg_28:readdata -> mm_interconnect_0:chrom_seg_28_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_28_s1_address;                // mm_interconnect_0:chrom_seg_28_s1_address -> chrom_seg_28:address
	wire         mm_interconnect_0_chrom_seg_28_s1_write;                  // mm_interconnect_0:chrom_seg_28_s1_write -> chrom_seg_28:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_28_s1_writedata;              // mm_interconnect_0:chrom_seg_28_s1_writedata -> chrom_seg_28:writedata
	wire         mm_interconnect_0_chrom_seg_29_s1_chipselect;             // mm_interconnect_0:chrom_seg_29_s1_chipselect -> chrom_seg_29:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_29_s1_readdata;               // chrom_seg_29:readdata -> mm_interconnect_0:chrom_seg_29_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_29_s1_address;                // mm_interconnect_0:chrom_seg_29_s1_address -> chrom_seg_29:address
	wire         mm_interconnect_0_chrom_seg_29_s1_write;                  // mm_interconnect_0:chrom_seg_29_s1_write -> chrom_seg_29:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_29_s1_writedata;              // mm_interconnect_0:chrom_seg_29_s1_writedata -> chrom_seg_29:writedata
	wire         mm_interconnect_0_chrom_seg_30_s1_chipselect;             // mm_interconnect_0:chrom_seg_30_s1_chipselect -> chrom_seg_30:chipselect
	wire  [31:0] mm_interconnect_0_chrom_seg_30_s1_readdata;               // chrom_seg_30:readdata -> mm_interconnect_0:chrom_seg_30_s1_readdata
	wire   [1:0] mm_interconnect_0_chrom_seg_30_s1_address;                // mm_interconnect_0:chrom_seg_30_s1_address -> chrom_seg_30:address
	wire         mm_interconnect_0_chrom_seg_30_s1_write;                  // mm_interconnect_0:chrom_seg_30_s1_write -> chrom_seg_30:write_n
	wire  [31:0] mm_interconnect_0_chrom_seg_30_s1_writedata;              // mm_interconnect_0:chrom_seg_30_s1_writedata -> chrom_seg_30:writedata
	wire         mm_interconnect_0_start_processing_chrom_s1_chipselect;   // mm_interconnect_0:start_processing_chrom_s1_chipselect -> start_processing_chrom:chipselect
	wire  [31:0] mm_interconnect_0_start_processing_chrom_s1_readdata;     // start_processing_chrom:readdata -> mm_interconnect_0:start_processing_chrom_s1_readdata
	wire   [1:0] mm_interconnect_0_start_processing_chrom_s1_address;      // mm_interconnect_0:start_processing_chrom_s1_address -> start_processing_chrom:address
	wire         mm_interconnect_0_start_processing_chrom_s1_write;        // mm_interconnect_0:start_processing_chrom_s1_write -> start_processing_chrom:write_n
	wire  [31:0] mm_interconnect_0_start_processing_chrom_s1_writedata;    // mm_interconnect_0:start_processing_chrom_s1_writedata -> start_processing_chrom:writedata
	wire  [31:0] mm_interconnect_0_done_processing_chrom_s1_readdata;      // done_processing_chrom:readdata -> mm_interconnect_0:done_processing_chrom_s1_readdata
	wire   [1:0] mm_interconnect_0_done_processing_chrom_s1_address;       // mm_interconnect_0:done_processing_chrom_s1_address -> done_processing_chrom:address
	wire  [31:0] mm_interconnect_0_ready_to_process_s1_readdata;           // ready_to_process:readdata -> mm_interconnect_0:ready_to_process_s1_readdata
	wire   [1:0] mm_interconnect_0_ready_to_process_s1_address;            // mm_interconnect_0:ready_to_process_s1_address -> ready_to_process:address
	wire         mm_interconnect_0_done_processing_feedback_s1_chipselect; // mm_interconnect_0:done_processing_feedback_s1_chipselect -> done_processing_feedback:chipselect
	wire  [31:0] mm_interconnect_0_done_processing_feedback_s1_readdata;   // done_processing_feedback:readdata -> mm_interconnect_0:done_processing_feedback_s1_readdata
	wire   [1:0] mm_interconnect_0_done_processing_feedback_s1_address;    // mm_interconnect_0:done_processing_feedback_s1_address -> done_processing_feedback:address
	wire         mm_interconnect_0_done_processing_feedback_s1_write;      // mm_interconnect_0:done_processing_feedback_s1_write -> done_processing_feedback:write_n
	wire  [31:0] mm_interconnect_0_done_processing_feedback_s1_writedata;  // mm_interconnect_0:done_processing_feedback_s1_writedata -> done_processing_feedback:writedata
	wire  [31:0] mm_interconnect_0_error_sum_0_s1_readdata;                // error_sum_0:readdata -> mm_interconnect_0:error_sum_0_s1_readdata
	wire   [1:0] mm_interconnect_0_error_sum_0_s1_address;                 // mm_interconnect_0:error_sum_0_s1_address -> error_sum_0:address
	wire  [31:0] mm_interconnect_0_error_sum_1_s1_readdata;                // error_sum_1:readdata -> mm_interconnect_0:error_sum_1_s1_readdata
	wire   [1:0] mm_interconnect_0_error_sum_1_s1_address;                 // mm_interconnect_0:error_sum_1_s1_address -> error_sum_1:address
	wire  [31:0] mm_interconnect_0_error_sum_2_s1_readdata;                // error_sum_2:readdata -> mm_interconnect_0:error_sum_2_s1_readdata
	wire   [1:0] mm_interconnect_0_error_sum_2_s1_address;                 // mm_interconnect_0:error_sum_2_s1_address -> error_sum_2:address
	wire  [31:0] mm_interconnect_0_error_sum_3_s1_readdata;                // error_sum_3:readdata -> mm_interconnect_0:error_sum_3_s1_readdata
	wire   [1:0] mm_interconnect_0_error_sum_3_s1_address;                 // mm_interconnect_0:error_sum_3_s1_address -> error_sum_3:address
	wire  [31:0] mm_interconnect_0_error_sum_4_s1_readdata;                // error_sum_4:readdata -> mm_interconnect_0:error_sum_4_s1_readdata
	wire   [1:0] mm_interconnect_0_error_sum_4_s1_address;                 // mm_interconnect_0:error_sum_4_s1_address -> error_sum_4:address
	wire  [31:0] mm_interconnect_0_error_sum_5_s1_readdata;                // error_sum_5:readdata -> mm_interconnect_0:error_sum_5_s1_readdata
	wire   [1:0] mm_interconnect_0_error_sum_5_s1_address;                 // mm_interconnect_0:error_sum_5_s1_address -> error_sum_5:address
	wire  [31:0] mm_interconnect_0_error_sum_6_s1_readdata;                // error_sum_6:readdata -> mm_interconnect_0:error_sum_6_s1_readdata
	wire   [1:0] mm_interconnect_0_error_sum_6_s1_address;                 // mm_interconnect_0:error_sum_6_s1_address -> error_sum_6:address
	wire  [31:0] mm_interconnect_0_error_sum_7_s1_readdata;                // error_sum_7:readdata -> mm_interconnect_0:error_sum_7_s1_readdata
	wire   [1:0] mm_interconnect_0_error_sum_7_s1_address;                 // mm_interconnect_0:error_sum_7_s1_address -> error_sum_7:address
	wire         mm_interconnect_0_input_sequence_0_s1_chipselect;         // mm_interconnect_0:input_sequence_0_s1_chipselect -> input_sequence_0:chipselect
	wire  [31:0] mm_interconnect_0_input_sequence_0_s1_readdata;           // input_sequence_0:readdata -> mm_interconnect_0:input_sequence_0_s1_readdata
	wire   [1:0] mm_interconnect_0_input_sequence_0_s1_address;            // mm_interconnect_0:input_sequence_0_s1_address -> input_sequence_0:address
	wire         mm_interconnect_0_input_sequence_0_s1_write;              // mm_interconnect_0:input_sequence_0_s1_write -> input_sequence_0:write_n
	wire  [31:0] mm_interconnect_0_input_sequence_0_s1_writedata;          // mm_interconnect_0:input_sequence_0_s1_writedata -> input_sequence_0:writedata
	wire         mm_interconnect_0_valid_output_0_s1_chipselect;           // mm_interconnect_0:valid_output_0_s1_chipselect -> valid_output_0:chipselect
	wire  [31:0] mm_interconnect_0_valid_output_0_s1_readdata;             // valid_output_0:readdata -> mm_interconnect_0:valid_output_0_s1_readdata
	wire   [1:0] mm_interconnect_0_valid_output_0_s1_address;              // mm_interconnect_0:valid_output_0_s1_address -> valid_output_0:address
	wire         mm_interconnect_0_valid_output_0_s1_write;                // mm_interconnect_0:valid_output_0_s1_write -> valid_output_0:write_n
	wire  [31:0] mm_interconnect_0_valid_output_0_s1_writedata;            // mm_interconnect_0:valid_output_0_s1_writedata -> valid_output_0:writedata
	wire         mm_interconnect_0_sequences_to_process_s1_chipselect;     // mm_interconnect_0:sequences_to_process_s1_chipselect -> sequences_to_process:chipselect
	wire  [31:0] mm_interconnect_0_sequences_to_process_s1_readdata;       // sequences_to_process:readdata -> mm_interconnect_0:sequences_to_process_s1_readdata
	wire   [1:0] mm_interconnect_0_sequences_to_process_s1_address;        // mm_interconnect_0:sequences_to_process_s1_address -> sequences_to_process:address
	wire         mm_interconnect_0_sequences_to_process_s1_write;          // mm_interconnect_0:sequences_to_process_s1_write -> sequences_to_process:write_n
	wire  [31:0] mm_interconnect_0_sequences_to_process_s1_writedata;      // mm_interconnect_0:sequences_to_process_s1_writedata -> sequences_to_process:writedata
	wire         mm_interconnect_0_two_port_mem_s1_chipselect;             // mm_interconnect_0:two_port_mem_s1_chipselect -> two_port_mem:chipselect
	wire  [31:0] mm_interconnect_0_two_port_mem_s1_readdata;               // two_port_mem:readdata -> mm_interconnect_0:two_port_mem_s1_readdata
	wire  [14:0] mm_interconnect_0_two_port_mem_s1_address;                // mm_interconnect_0:two_port_mem_s1_address -> two_port_mem:address
	wire   [3:0] mm_interconnect_0_two_port_mem_s1_byteenable;             // mm_interconnect_0:two_port_mem_s1_byteenable -> two_port_mem:byteenable
	wire         mm_interconnect_0_two_port_mem_s1_write;                  // mm_interconnect_0:two_port_mem_s1_write -> two_port_mem:write
	wire  [31:0] mm_interconnect_0_two_port_mem_s1_writedata;              // mm_interconnect_0:two_port_mem_s1_writedata -> two_port_mem:writedata
	wire         mm_interconnect_0_two_port_mem_s1_clken;                  // mm_interconnect_0:two_port_mem_s1_clken -> two_port_mem:clken
	wire         mm_interconnect_0_two_port_mem_correct_s1_chipselect;     // mm_interconnect_0:two_port_mem_correct_s1_chipselect -> two_port_mem_correct:chipselect
	wire  [31:0] mm_interconnect_0_two_port_mem_correct_s1_readdata;       // two_port_mem_correct:readdata -> mm_interconnect_0:two_port_mem_correct_s1_readdata
	wire  [14:0] mm_interconnect_0_two_port_mem_correct_s1_address;        // mm_interconnect_0:two_port_mem_correct_s1_address -> two_port_mem_correct:address
	wire   [3:0] mm_interconnect_0_two_port_mem_correct_s1_byteenable;     // mm_interconnect_0:two_port_mem_correct_s1_byteenable -> two_port_mem_correct:byteenable
	wire         mm_interconnect_0_two_port_mem_correct_s1_write;          // mm_interconnect_0:two_port_mem_correct_s1_write -> two_port_mem_correct:write
	wire  [31:0] mm_interconnect_0_two_port_mem_correct_s1_writedata;      // mm_interconnect_0:two_port_mem_correct_s1_writedata -> two_port_mem_correct:writedata
	wire         mm_interconnect_0_two_port_mem_correct_s1_clken;          // mm_interconnect_0:two_port_mem_correct_s1_clken -> two_port_mem_correct:clken
	wire         mm_interconnect_0_expected_output_0_s1_chipselect;        // mm_interconnect_0:expected_output_0_s1_chipselect -> expected_output_0:chipselect
	wire  [31:0] mm_interconnect_0_expected_output_0_s1_readdata;          // expected_output_0:readdata -> mm_interconnect_0:expected_output_0_s1_readdata
	wire   [1:0] mm_interconnect_0_expected_output_0_s1_address;           // mm_interconnect_0:expected_output_0_s1_address -> expected_output_0:address
	wire         mm_interconnect_0_expected_output_0_s1_write;             // mm_interconnect_0:expected_output_0_s1_write -> expected_output_0:write_n
	wire  [31:0] mm_interconnect_0_expected_output_0_s1_writedata;         // mm_interconnect_0:expected_output_0_s1_writedata -> expected_output_0:writedata
	wire         mm_interconnect_0_writesample_s1_chipselect;              // mm_interconnect_0:writeSample_s1_chipselect -> writeSample:chipselect
	wire  [31:0] mm_interconnect_0_writesample_s1_readdata;                // writeSample:readdata -> mm_interconnect_0:writeSample_s1_readdata
	wire   [1:0] mm_interconnect_0_writesample_s1_address;                 // mm_interconnect_0:writeSample_s1_address -> writeSample:address
	wire         mm_interconnect_0_writesample_s1_write;                   // mm_interconnect_0:writeSample_s1_write -> writeSample:write_n
	wire  [31:0] mm_interconnect_0_writesample_s1_writedata;               // mm_interconnect_0:writeSample_s1_writedata -> writeSample:writedata
	wire         mm_interconnect_0_sampleindex_s1_chipselect;              // mm_interconnect_0:sampleIndex_s1_chipselect -> sampleIndex:chipselect
	wire  [31:0] mm_interconnect_0_sampleindex_s1_readdata;                // sampleIndex:readdata -> mm_interconnect_0:sampleIndex_s1_readdata
	wire   [1:0] mm_interconnect_0_sampleindex_s1_address;                 // mm_interconnect_0:sampleIndex_s1_address -> sampleIndex:address
	wire         mm_interconnect_0_sampleindex_s1_write;                   // mm_interconnect_0:sampleIndex_s1_write -> sampleIndex:write_n
	wire  [31:0] mm_interconnect_0_sampleindex_s1_writedata;               // mm_interconnect_0:sampleIndex_s1_writedata -> sampleIndex:writedata
	wire  [31:0] mm_interconnect_0_nextsample_s1_readdata;                 // nextSample:readdata -> mm_interconnect_0:nextSample_s1_readdata
	wire   [1:0] mm_interconnect_0_nextsample_s1_address;                  // mm_interconnect_0:nextSample_s1_address -> nextSample:address
	wire         mm_interconnect_0_preparingnextsample_s1_chipselect;      // mm_interconnect_0:preparingNextSample_s1_chipselect -> preparingNextSample:chipselect
	wire  [31:0] mm_interconnect_0_preparingnextsample_s1_readdata;        // preparingNextSample:readdata -> mm_interconnect_0:preparingNextSample_s1_readdata
	wire   [1:0] mm_interconnect_0_preparingnextsample_s1_address;         // mm_interconnect_0:preparingNextSample_s1_address -> preparingNextSample:address
	wire         mm_interconnect_0_preparingnextsample_s1_write;           // mm_interconnect_0:preparingNextSample_s1_write -> preparingNextSample:write_n
	wire  [31:0] mm_interconnect_0_preparingnextsample_s1_writedata;       // mm_interconnect_0:preparingNextSample_s1_writedata -> preparingNextSample:writedata
	wire         rst_controller_reset_out_reset;                           // rst_controller:reset_out -> [chrom_seg_0:reset_n, chrom_seg_10:reset_n, chrom_seg_11:reset_n, chrom_seg_12:reset_n, chrom_seg_13:reset_n, chrom_seg_14:reset_n, chrom_seg_15:reset_n, chrom_seg_16:reset_n, chrom_seg_17:reset_n, chrom_seg_18:reset_n, chrom_seg_19:reset_n, chrom_seg_1:reset_n, chrom_seg_20:reset_n, chrom_seg_21:reset_n, chrom_seg_22:reset_n, chrom_seg_23:reset_n, chrom_seg_24:reset_n, chrom_seg_25:reset_n, chrom_seg_26:reset_n, chrom_seg_27:reset_n, chrom_seg_28:reset_n, chrom_seg_29:reset_n, chrom_seg_2:reset_n, chrom_seg_30:reset_n, chrom_seg_3:reset_n, chrom_seg_4:reset_n, chrom_seg_5:reset_n, chrom_seg_6:reset_n, chrom_seg_7:reset_n, chrom_seg_8:reset_n, chrom_seg_9:reset_n, done_processing_chrom:reset_n, done_processing_feedback:reset_n, error_sum_0:reset_n, error_sum_1:reset_n, error_sum_2:reset_n, error_sum_3:reset_n, error_sum_4:reset_n, error_sum_5:reset_n, error_sum_6:reset_n, error_sum_7:reset_n, expected_output_0:reset_n, input_sequence_0:reset_n, mm_interconnect_0:chrom_seg_0_reset_reset_bridge_in_reset_reset, nextSample:reset_n, preparingNextSample:reset_n, ready_to_process:reset_n, rst_translator:in_reset, sampleIndex:reset_n, sequences_to_process:reset_n, start_processing_chrom:reset_n, two_port_mem:reset, two_port_mem:reset2, two_port_mem_correct:reset, two_port_mem_correct:reset2, valid_output_0:reset_n, writeSample:reset_n]
	wire         rst_controller_reset_out_reset_req;                       // rst_controller:reset_req -> [rst_translator:reset_req_in, two_port_mem:reset_req, two_port_mem:reset_req2, two_port_mem_correct:reset_req, two_port_mem_correct:reset_req2]
	wire         hps_0_h2f_reset_reset;                                    // hps_0:h2f_rst_n -> rst_controller:reset_in0

	testeio_chrom_seg_0 chrom_seg_0 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_0_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_0_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_1 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_1_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_1_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_10 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_10_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_10_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_10_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_10_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_10_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_10_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_11 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_11_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_11_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_11_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_11_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_11_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_11_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_12 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_12_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_12_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_12_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_12_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_12_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_12_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_13 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_13_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_13_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_13_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_13_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_13_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_13_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_14 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_14_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_14_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_14_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_14_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_14_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_14_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_15 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_15_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_15_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_15_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_15_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_15_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_15_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_16 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_16_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_16_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_16_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_16_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_16_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_16_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_17 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_17_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_17_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_17_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_17_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_17_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_17_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_18 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_18_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_18_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_18_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_18_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_18_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_18_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_19 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_19_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_19_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_19_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_19_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_19_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_19_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_2 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_2_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_2_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_20 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_20_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_20_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_20_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_20_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_20_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_20_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_21 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_21_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_21_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_21_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_21_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_21_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_21_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_22 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_22_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_22_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_22_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_22_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_22_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_22_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_23 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_23_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_23_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_23_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_23_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_23_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_23_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_24 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_24_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_24_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_24_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_24_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_24_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_24_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_25 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_25_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_25_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_25_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_25_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_25_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_25_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_26 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_26_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_26_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_26_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_26_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_26_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_26_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_27 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_27_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_27_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_27_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_27_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_27_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_27_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_28 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_28_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_28_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_28_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_28_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_28_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_28_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_29 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_29_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_29_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_29_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_29_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_29_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_29_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_3 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_3_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_3_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_30 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_30_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_30_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_30_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_30_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_30_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_30_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_4 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_4_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_4_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_5 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_5_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_5_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_6 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_6_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_6_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_7 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_7_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_7_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_8 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_8_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_8_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 chrom_seg_9 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_chrom_seg_9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chrom_seg_9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chrom_seg_9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chrom_seg_9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chrom_seg_9_s1_readdata),   //                    .readdata
		.out_port   (chrom_seg_9_export)                           // external_connection.export
	);

	testeio_done_processing_chrom done_processing_chrom (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address  (mm_interconnect_0_done_processing_chrom_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_done_processing_chrom_s1_readdata), //                    .readdata
		.in_port  (done_processing_chrom_export)                         // external_connection.export
	);

	testeio_done_processing_feedback done_processing_feedback (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                          //               reset.reset_n
		.address    (mm_interconnect_0_done_processing_feedback_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_done_processing_feedback_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_done_processing_feedback_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_done_processing_feedback_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_done_processing_feedback_s1_readdata),   //                    .readdata
		.out_port   (done_processing_feedback_export)                           // external_connection.export
	);

	testeio_error_sum_0 error_sum_0 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_error_sum_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_error_sum_0_s1_readdata), //                    .readdata
		.in_port  (error_sum_0_export)                         // external_connection.export
	);

	testeio_error_sum_0 error_sum_1 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_error_sum_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_error_sum_1_s1_readdata), //                    .readdata
		.in_port  (error_sum_1_export)                         // external_connection.export
	);

	testeio_error_sum_0 error_sum_2 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_error_sum_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_error_sum_2_s1_readdata), //                    .readdata
		.in_port  (error_sum_2_export)                         // external_connection.export
	);

	testeio_error_sum_0 error_sum_3 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_error_sum_3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_error_sum_3_s1_readdata), //                    .readdata
		.in_port  (error_sum_3_export)                         // external_connection.export
	);

	testeio_error_sum_0 error_sum_4 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_error_sum_4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_error_sum_4_s1_readdata), //                    .readdata
		.in_port  (error_sum_4_export)                         // external_connection.export
	);

	testeio_error_sum_0 error_sum_5 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_error_sum_5_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_error_sum_5_s1_readdata), //                    .readdata
		.in_port  (error_sum_5_export)                         // external_connection.export
	);

	testeio_error_sum_0 error_sum_6 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_error_sum_6_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_error_sum_6_s1_readdata), //                    .readdata
		.in_port  (error_sum_6_export)                         // external_connection.export
	);

	testeio_error_sum_0 error_sum_7 (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_error_sum_7_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_error_sum_7_s1_readdata), //                    .readdata
		.in_port  (error_sum_7_export)                         // external_connection.export
	);

	testeio_chrom_seg_0 expected_output_0 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_expected_output_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_expected_output_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_expected_output_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_expected_output_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_expected_output_0_s1_readdata),   //                    .readdata
		.out_port   (expected_output_0_export)                           // external_connection.export
	);

	testeio_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.mem_a                    (memory_mem_a),                    //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                   //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                   //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                  //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),              //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                   //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                  //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                   //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK), //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL), //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL), //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK), //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),   //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),     //                  .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),     //                  .hps_io_uart0_inst_TX
		.h2f_rst_n                (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                         //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                //                  .awaddr
		.h2f_AWLEN                (),                                //                  .awlen
		.h2f_AWSIZE               (),                                //                  .awsize
		.h2f_AWBURST              (),                                //                  .awburst
		.h2f_AWLOCK               (),                                //                  .awlock
		.h2f_AWCACHE              (),                                //                  .awcache
		.h2f_AWPROT               (),                                //                  .awprot
		.h2f_AWVALID              (),                                //                  .awvalid
		.h2f_AWREADY              (),                                //                  .awready
		.h2f_WID                  (),                                //                  .wid
		.h2f_WDATA                (),                                //                  .wdata
		.h2f_WSTRB                (),                                //                  .wstrb
		.h2f_WLAST                (),                                //                  .wlast
		.h2f_WVALID               (),                                //                  .wvalid
		.h2f_WREADY               (),                                //                  .wready
		.h2f_BID                  (),                                //                  .bid
		.h2f_BRESP                (),                                //                  .bresp
		.h2f_BVALID               (),                                //                  .bvalid
		.h2f_BREADY               (),                                //                  .bready
		.h2f_ARID                 (),                                //                  .arid
		.h2f_ARADDR               (),                                //                  .araddr
		.h2f_ARLEN                (),                                //                  .arlen
		.h2f_ARSIZE               (),                                //                  .arsize
		.h2f_ARBURST              (),                                //                  .arburst
		.h2f_ARLOCK               (),                                //                  .arlock
		.h2f_ARCACHE              (),                                //                  .arcache
		.h2f_ARPROT               (),                                //                  .arprot
		.h2f_ARVALID              (),                                //                  .arvalid
		.h2f_ARREADY              (),                                //                  .arready
		.h2f_RID                  (),                                //                  .rid
		.h2f_RDATA                (),                                //                  .rdata
		.h2f_RRESP                (),                                //                  .rresp
		.h2f_RLAST                (),                                //                  .rlast
		.h2f_RVALID               (),                                //                  .rvalid
		.h2f_RREADY               (),                                //                  .rready
		.f2h_axi_clk              (clk_clk),                         //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                //                  .awaddr
		.f2h_AWLEN                (),                                //                  .awlen
		.f2h_AWSIZE               (),                                //                  .awsize
		.f2h_AWBURST              (),                                //                  .awburst
		.f2h_AWLOCK               (),                                //                  .awlock
		.f2h_AWCACHE              (),                                //                  .awcache
		.f2h_AWPROT               (),                                //                  .awprot
		.f2h_AWVALID              (),                                //                  .awvalid
		.f2h_AWREADY              (),                                //                  .awready
		.f2h_AWUSER               (),                                //                  .awuser
		.f2h_WID                  (),                                //                  .wid
		.f2h_WDATA                (),                                //                  .wdata
		.f2h_WSTRB                (),                                //                  .wstrb
		.f2h_WLAST                (),                                //                  .wlast
		.f2h_WVALID               (),                                //                  .wvalid
		.f2h_WREADY               (),                                //                  .wready
		.f2h_BID                  (),                                //                  .bid
		.f2h_BRESP                (),                                //                  .bresp
		.f2h_BVALID               (),                                //                  .bvalid
		.f2h_BREADY               (),                                //                  .bready
		.f2h_ARID                 (),                                //                  .arid
		.f2h_ARADDR               (),                                //                  .araddr
		.f2h_ARLEN                (),                                //                  .arlen
		.f2h_ARSIZE               (),                                //                  .arsize
		.f2h_ARBURST              (),                                //                  .arburst
		.f2h_ARLOCK               (),                                //                  .arlock
		.f2h_ARCACHE              (),                                //                  .arcache
		.f2h_ARPROT               (),                                //                  .arprot
		.f2h_ARVALID              (),                                //                  .arvalid
		.f2h_ARREADY              (),                                //                  .arready
		.f2h_ARUSER               (),                                //                  .aruser
		.f2h_RID                  (),                                //                  .rid
		.f2h_RDATA                (),                                //                  .rdata
		.f2h_RRESP                (),                                //                  .rresp
		.f2h_RLAST                (),                                //                  .rlast
		.f2h_RVALID               (),                                //                  .rvalid
		.f2h_RREADY               (),                                //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                         //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready)   //                  .rready
	);

	testeio_chrom_seg_0 input_sequence_0 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_input_sequence_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_input_sequence_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_input_sequence_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_input_sequence_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_input_sequence_0_s1_readdata),   //                    .readdata
		.out_port   (input_sequence_0_export)                           // external_connection.export
	);

	testeio_error_sum_0 nextsample (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_nextsample_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_nextsample_s1_readdata), //                    .readdata
		.in_port  (nextsample_export)                         // external_connection.export
	);

	testeio_chrom_seg_0 preparingnextsample (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (mm_interconnect_0_preparingnextsample_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_preparingnextsample_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_preparingnextsample_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_preparingnextsample_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_preparingnextsample_s1_readdata),   //                    .readdata
		.out_port   (preparingnextsample_export)                           // external_connection.export
	);

	testeio_done_processing_chrom ready_to_process (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_ready_to_process_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ready_to_process_s1_readdata), //                    .readdata
		.in_port  (ready_to_process_export)                         // external_connection.export
	);

	testeio_chrom_seg_0 sampleindex (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_sampleindex_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sampleindex_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sampleindex_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sampleindex_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sampleindex_s1_readdata),   //                    .readdata
		.out_port   (sampleindex_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 sequences_to_process (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (mm_interconnect_0_sequences_to_process_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sequences_to_process_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sequences_to_process_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sequences_to_process_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sequences_to_process_s1_readdata),   //                    .readdata
		.out_port   (sequences_to_process_export)                           // external_connection.export
	);

	testeio_done_processing_feedback start_processing_chrom (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address    (mm_interconnect_0_start_processing_chrom_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_processing_chrom_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_processing_chrom_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_processing_chrom_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_processing_chrom_s1_readdata),   //                    .readdata
		.out_port   (start_processing_chrom_export)                           // external_connection.export
	);

	testeio_two_port_mem two_port_mem (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_two_port_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_two_port_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_two_port_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_two_port_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_0_two_port_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_two_port_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_two_port_mem_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),           //       .reset_req
		.address2    (mem_s2_address),                               //     s2.address
		.chipselect2 (mem_s2_chipselect),                            //       .chipselect
		.clken2      (mem_s2_clken),                                 //       .clken
		.write2      (mem_s2_write),                                 //       .write
		.readdata2   (mem_s2_readdata),                              //       .readdata
		.writedata2  (mem_s2_writedata),                             //       .writedata
		.byteenable2 (mem_s2_byteenable),                            //       .byteenable
		.clk2        (clk_clk),                                      //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),               // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                          // (terminated)
	);

	testeio_two_port_mem_correct two_port_mem_correct (
		.clk         (clk_clk),                                              //   clk1.clk
		.address     (mm_interconnect_0_two_port_mem_correct_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_two_port_mem_correct_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_two_port_mem_correct_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_two_port_mem_correct_s1_write),      //       .write
		.readdata    (mm_interconnect_0_two_port_mem_correct_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_two_port_mem_correct_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_two_port_mem_correct_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),                   //       .reset_req
		.address2    (correct_mem_s2_address),                               //     s2.address
		.chipselect2 (correct_mem_s2_chipselect),                            //       .chipselect
		.clken2      (correct_mem_s2_clken),                                 //       .clken
		.write2      (correct_mem_s2_write),                                 //       .write
		.readdata2   (correct_mem_s2_readdata),                              //       .readdata
		.writedata2  (correct_mem_s2_writedata),                             //       .writedata
		.byteenable2 (correct_mem_s2_byteenable),                            //       .byteenable
		.clk2        (clk_clk),                                              //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                       // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),                   //       .reset_req
		.freeze      (1'b0)                                                  // (terminated)
	);

	testeio_chrom_seg_0 valid_output_0 (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_valid_output_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_valid_output_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_valid_output_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_valid_output_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_valid_output_0_s1_readdata),   //                    .readdata
		.out_port   (valid_output_0_export)                           // external_connection.export
	);

	testeio_chrom_seg_0 writesample (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_writesample_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_writesample_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_writesample_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_writesample_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_writesample_s1_readdata),   //                    .readdata
		.out_port   (writesample_export)                           // external_connection.export
	);

	testeio_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                  (hps_0_h2f_lw_axi_master_awid),                             //                 hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                (hps_0_h2f_lw_axi_master_awaddr),                           //                                        .awaddr
		.hps_0_h2f_lw_axi_master_awlen                 (hps_0_h2f_lw_axi_master_awlen),                            //                                        .awlen
		.hps_0_h2f_lw_axi_master_awsize                (hps_0_h2f_lw_axi_master_awsize),                           //                                        .awsize
		.hps_0_h2f_lw_axi_master_awburst               (hps_0_h2f_lw_axi_master_awburst),                          //                                        .awburst
		.hps_0_h2f_lw_axi_master_awlock                (hps_0_h2f_lw_axi_master_awlock),                           //                                        .awlock
		.hps_0_h2f_lw_axi_master_awcache               (hps_0_h2f_lw_axi_master_awcache),                          //                                        .awcache
		.hps_0_h2f_lw_axi_master_awprot                (hps_0_h2f_lw_axi_master_awprot),                           //                                        .awprot
		.hps_0_h2f_lw_axi_master_awvalid               (hps_0_h2f_lw_axi_master_awvalid),                          //                                        .awvalid
		.hps_0_h2f_lw_axi_master_awready               (hps_0_h2f_lw_axi_master_awready),                          //                                        .awready
		.hps_0_h2f_lw_axi_master_wid                   (hps_0_h2f_lw_axi_master_wid),                              //                                        .wid
		.hps_0_h2f_lw_axi_master_wdata                 (hps_0_h2f_lw_axi_master_wdata),                            //                                        .wdata
		.hps_0_h2f_lw_axi_master_wstrb                 (hps_0_h2f_lw_axi_master_wstrb),                            //                                        .wstrb
		.hps_0_h2f_lw_axi_master_wlast                 (hps_0_h2f_lw_axi_master_wlast),                            //                                        .wlast
		.hps_0_h2f_lw_axi_master_wvalid                (hps_0_h2f_lw_axi_master_wvalid),                           //                                        .wvalid
		.hps_0_h2f_lw_axi_master_wready                (hps_0_h2f_lw_axi_master_wready),                           //                                        .wready
		.hps_0_h2f_lw_axi_master_bid                   (hps_0_h2f_lw_axi_master_bid),                              //                                        .bid
		.hps_0_h2f_lw_axi_master_bresp                 (hps_0_h2f_lw_axi_master_bresp),                            //                                        .bresp
		.hps_0_h2f_lw_axi_master_bvalid                (hps_0_h2f_lw_axi_master_bvalid),                           //                                        .bvalid
		.hps_0_h2f_lw_axi_master_bready                (hps_0_h2f_lw_axi_master_bready),                           //                                        .bready
		.hps_0_h2f_lw_axi_master_arid                  (hps_0_h2f_lw_axi_master_arid),                             //                                        .arid
		.hps_0_h2f_lw_axi_master_araddr                (hps_0_h2f_lw_axi_master_araddr),                           //                                        .araddr
		.hps_0_h2f_lw_axi_master_arlen                 (hps_0_h2f_lw_axi_master_arlen),                            //                                        .arlen
		.hps_0_h2f_lw_axi_master_arsize                (hps_0_h2f_lw_axi_master_arsize),                           //                                        .arsize
		.hps_0_h2f_lw_axi_master_arburst               (hps_0_h2f_lw_axi_master_arburst),                          //                                        .arburst
		.hps_0_h2f_lw_axi_master_arlock                (hps_0_h2f_lw_axi_master_arlock),                           //                                        .arlock
		.hps_0_h2f_lw_axi_master_arcache               (hps_0_h2f_lw_axi_master_arcache),                          //                                        .arcache
		.hps_0_h2f_lw_axi_master_arprot                (hps_0_h2f_lw_axi_master_arprot),                           //                                        .arprot
		.hps_0_h2f_lw_axi_master_arvalid               (hps_0_h2f_lw_axi_master_arvalid),                          //                                        .arvalid
		.hps_0_h2f_lw_axi_master_arready               (hps_0_h2f_lw_axi_master_arready),                          //                                        .arready
		.hps_0_h2f_lw_axi_master_rid                   (hps_0_h2f_lw_axi_master_rid),                              //                                        .rid
		.hps_0_h2f_lw_axi_master_rdata                 (hps_0_h2f_lw_axi_master_rdata),                            //                                        .rdata
		.hps_0_h2f_lw_axi_master_rresp                 (hps_0_h2f_lw_axi_master_rresp),                            //                                        .rresp
		.hps_0_h2f_lw_axi_master_rlast                 (hps_0_h2f_lw_axi_master_rlast),                            //                                        .rlast
		.hps_0_h2f_lw_axi_master_rvalid                (hps_0_h2f_lw_axi_master_rvalid),                           //                                        .rvalid
		.hps_0_h2f_lw_axi_master_rready                (hps_0_h2f_lw_axi_master_rready),                           //                                        .rready
		.clk_0_clk_clk                                 (clk_clk),                                                  //                               clk_0_clk.clk
		.chrom_seg_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                           // chrom_seg_0_reset_reset_bridge_in_reset.reset
		.chrom_seg_0_s1_address                        (mm_interconnect_0_chrom_seg_0_s1_address),                 //                          chrom_seg_0_s1.address
		.chrom_seg_0_s1_write                          (mm_interconnect_0_chrom_seg_0_s1_write),                   //                                        .write
		.chrom_seg_0_s1_readdata                       (mm_interconnect_0_chrom_seg_0_s1_readdata),                //                                        .readdata
		.chrom_seg_0_s1_writedata                      (mm_interconnect_0_chrom_seg_0_s1_writedata),               //                                        .writedata
		.chrom_seg_0_s1_chipselect                     (mm_interconnect_0_chrom_seg_0_s1_chipselect),              //                                        .chipselect
		.chrom_seg_1_s1_address                        (mm_interconnect_0_chrom_seg_1_s1_address),                 //                          chrom_seg_1_s1.address
		.chrom_seg_1_s1_write                          (mm_interconnect_0_chrom_seg_1_s1_write),                   //                                        .write
		.chrom_seg_1_s1_readdata                       (mm_interconnect_0_chrom_seg_1_s1_readdata),                //                                        .readdata
		.chrom_seg_1_s1_writedata                      (mm_interconnect_0_chrom_seg_1_s1_writedata),               //                                        .writedata
		.chrom_seg_1_s1_chipselect                     (mm_interconnect_0_chrom_seg_1_s1_chipselect),              //                                        .chipselect
		.chrom_seg_10_s1_address                       (mm_interconnect_0_chrom_seg_10_s1_address),                //                         chrom_seg_10_s1.address
		.chrom_seg_10_s1_write                         (mm_interconnect_0_chrom_seg_10_s1_write),                  //                                        .write
		.chrom_seg_10_s1_readdata                      (mm_interconnect_0_chrom_seg_10_s1_readdata),               //                                        .readdata
		.chrom_seg_10_s1_writedata                     (mm_interconnect_0_chrom_seg_10_s1_writedata),              //                                        .writedata
		.chrom_seg_10_s1_chipselect                    (mm_interconnect_0_chrom_seg_10_s1_chipselect),             //                                        .chipselect
		.chrom_seg_11_s1_address                       (mm_interconnect_0_chrom_seg_11_s1_address),                //                         chrom_seg_11_s1.address
		.chrom_seg_11_s1_write                         (mm_interconnect_0_chrom_seg_11_s1_write),                  //                                        .write
		.chrom_seg_11_s1_readdata                      (mm_interconnect_0_chrom_seg_11_s1_readdata),               //                                        .readdata
		.chrom_seg_11_s1_writedata                     (mm_interconnect_0_chrom_seg_11_s1_writedata),              //                                        .writedata
		.chrom_seg_11_s1_chipselect                    (mm_interconnect_0_chrom_seg_11_s1_chipselect),             //                                        .chipselect
		.chrom_seg_12_s1_address                       (mm_interconnect_0_chrom_seg_12_s1_address),                //                         chrom_seg_12_s1.address
		.chrom_seg_12_s1_write                         (mm_interconnect_0_chrom_seg_12_s1_write),                  //                                        .write
		.chrom_seg_12_s1_readdata                      (mm_interconnect_0_chrom_seg_12_s1_readdata),               //                                        .readdata
		.chrom_seg_12_s1_writedata                     (mm_interconnect_0_chrom_seg_12_s1_writedata),              //                                        .writedata
		.chrom_seg_12_s1_chipselect                    (mm_interconnect_0_chrom_seg_12_s1_chipselect),             //                                        .chipselect
		.chrom_seg_13_s1_address                       (mm_interconnect_0_chrom_seg_13_s1_address),                //                         chrom_seg_13_s1.address
		.chrom_seg_13_s1_write                         (mm_interconnect_0_chrom_seg_13_s1_write),                  //                                        .write
		.chrom_seg_13_s1_readdata                      (mm_interconnect_0_chrom_seg_13_s1_readdata),               //                                        .readdata
		.chrom_seg_13_s1_writedata                     (mm_interconnect_0_chrom_seg_13_s1_writedata),              //                                        .writedata
		.chrom_seg_13_s1_chipselect                    (mm_interconnect_0_chrom_seg_13_s1_chipselect),             //                                        .chipselect
		.chrom_seg_14_s1_address                       (mm_interconnect_0_chrom_seg_14_s1_address),                //                         chrom_seg_14_s1.address
		.chrom_seg_14_s1_write                         (mm_interconnect_0_chrom_seg_14_s1_write),                  //                                        .write
		.chrom_seg_14_s1_readdata                      (mm_interconnect_0_chrom_seg_14_s1_readdata),               //                                        .readdata
		.chrom_seg_14_s1_writedata                     (mm_interconnect_0_chrom_seg_14_s1_writedata),              //                                        .writedata
		.chrom_seg_14_s1_chipselect                    (mm_interconnect_0_chrom_seg_14_s1_chipselect),             //                                        .chipselect
		.chrom_seg_15_s1_address                       (mm_interconnect_0_chrom_seg_15_s1_address),                //                         chrom_seg_15_s1.address
		.chrom_seg_15_s1_write                         (mm_interconnect_0_chrom_seg_15_s1_write),                  //                                        .write
		.chrom_seg_15_s1_readdata                      (mm_interconnect_0_chrom_seg_15_s1_readdata),               //                                        .readdata
		.chrom_seg_15_s1_writedata                     (mm_interconnect_0_chrom_seg_15_s1_writedata),              //                                        .writedata
		.chrom_seg_15_s1_chipselect                    (mm_interconnect_0_chrom_seg_15_s1_chipselect),             //                                        .chipselect
		.chrom_seg_16_s1_address                       (mm_interconnect_0_chrom_seg_16_s1_address),                //                         chrom_seg_16_s1.address
		.chrom_seg_16_s1_write                         (mm_interconnect_0_chrom_seg_16_s1_write),                  //                                        .write
		.chrom_seg_16_s1_readdata                      (mm_interconnect_0_chrom_seg_16_s1_readdata),               //                                        .readdata
		.chrom_seg_16_s1_writedata                     (mm_interconnect_0_chrom_seg_16_s1_writedata),              //                                        .writedata
		.chrom_seg_16_s1_chipselect                    (mm_interconnect_0_chrom_seg_16_s1_chipselect),             //                                        .chipselect
		.chrom_seg_17_s1_address                       (mm_interconnect_0_chrom_seg_17_s1_address),                //                         chrom_seg_17_s1.address
		.chrom_seg_17_s1_write                         (mm_interconnect_0_chrom_seg_17_s1_write),                  //                                        .write
		.chrom_seg_17_s1_readdata                      (mm_interconnect_0_chrom_seg_17_s1_readdata),               //                                        .readdata
		.chrom_seg_17_s1_writedata                     (mm_interconnect_0_chrom_seg_17_s1_writedata),              //                                        .writedata
		.chrom_seg_17_s1_chipselect                    (mm_interconnect_0_chrom_seg_17_s1_chipselect),             //                                        .chipselect
		.chrom_seg_18_s1_address                       (mm_interconnect_0_chrom_seg_18_s1_address),                //                         chrom_seg_18_s1.address
		.chrom_seg_18_s1_write                         (mm_interconnect_0_chrom_seg_18_s1_write),                  //                                        .write
		.chrom_seg_18_s1_readdata                      (mm_interconnect_0_chrom_seg_18_s1_readdata),               //                                        .readdata
		.chrom_seg_18_s1_writedata                     (mm_interconnect_0_chrom_seg_18_s1_writedata),              //                                        .writedata
		.chrom_seg_18_s1_chipselect                    (mm_interconnect_0_chrom_seg_18_s1_chipselect),             //                                        .chipselect
		.chrom_seg_19_s1_address                       (mm_interconnect_0_chrom_seg_19_s1_address),                //                         chrom_seg_19_s1.address
		.chrom_seg_19_s1_write                         (mm_interconnect_0_chrom_seg_19_s1_write),                  //                                        .write
		.chrom_seg_19_s1_readdata                      (mm_interconnect_0_chrom_seg_19_s1_readdata),               //                                        .readdata
		.chrom_seg_19_s1_writedata                     (mm_interconnect_0_chrom_seg_19_s1_writedata),              //                                        .writedata
		.chrom_seg_19_s1_chipselect                    (mm_interconnect_0_chrom_seg_19_s1_chipselect),             //                                        .chipselect
		.chrom_seg_2_s1_address                        (mm_interconnect_0_chrom_seg_2_s1_address),                 //                          chrom_seg_2_s1.address
		.chrom_seg_2_s1_write                          (mm_interconnect_0_chrom_seg_2_s1_write),                   //                                        .write
		.chrom_seg_2_s1_readdata                       (mm_interconnect_0_chrom_seg_2_s1_readdata),                //                                        .readdata
		.chrom_seg_2_s1_writedata                      (mm_interconnect_0_chrom_seg_2_s1_writedata),               //                                        .writedata
		.chrom_seg_2_s1_chipselect                     (mm_interconnect_0_chrom_seg_2_s1_chipselect),              //                                        .chipselect
		.chrom_seg_20_s1_address                       (mm_interconnect_0_chrom_seg_20_s1_address),                //                         chrom_seg_20_s1.address
		.chrom_seg_20_s1_write                         (mm_interconnect_0_chrom_seg_20_s1_write),                  //                                        .write
		.chrom_seg_20_s1_readdata                      (mm_interconnect_0_chrom_seg_20_s1_readdata),               //                                        .readdata
		.chrom_seg_20_s1_writedata                     (mm_interconnect_0_chrom_seg_20_s1_writedata),              //                                        .writedata
		.chrom_seg_20_s1_chipselect                    (mm_interconnect_0_chrom_seg_20_s1_chipselect),             //                                        .chipselect
		.chrom_seg_21_s1_address                       (mm_interconnect_0_chrom_seg_21_s1_address),                //                         chrom_seg_21_s1.address
		.chrom_seg_21_s1_write                         (mm_interconnect_0_chrom_seg_21_s1_write),                  //                                        .write
		.chrom_seg_21_s1_readdata                      (mm_interconnect_0_chrom_seg_21_s1_readdata),               //                                        .readdata
		.chrom_seg_21_s1_writedata                     (mm_interconnect_0_chrom_seg_21_s1_writedata),              //                                        .writedata
		.chrom_seg_21_s1_chipselect                    (mm_interconnect_0_chrom_seg_21_s1_chipselect),             //                                        .chipselect
		.chrom_seg_22_s1_address                       (mm_interconnect_0_chrom_seg_22_s1_address),                //                         chrom_seg_22_s1.address
		.chrom_seg_22_s1_write                         (mm_interconnect_0_chrom_seg_22_s1_write),                  //                                        .write
		.chrom_seg_22_s1_readdata                      (mm_interconnect_0_chrom_seg_22_s1_readdata),               //                                        .readdata
		.chrom_seg_22_s1_writedata                     (mm_interconnect_0_chrom_seg_22_s1_writedata),              //                                        .writedata
		.chrom_seg_22_s1_chipselect                    (mm_interconnect_0_chrom_seg_22_s1_chipselect),             //                                        .chipselect
		.chrom_seg_23_s1_address                       (mm_interconnect_0_chrom_seg_23_s1_address),                //                         chrom_seg_23_s1.address
		.chrom_seg_23_s1_write                         (mm_interconnect_0_chrom_seg_23_s1_write),                  //                                        .write
		.chrom_seg_23_s1_readdata                      (mm_interconnect_0_chrom_seg_23_s1_readdata),               //                                        .readdata
		.chrom_seg_23_s1_writedata                     (mm_interconnect_0_chrom_seg_23_s1_writedata),              //                                        .writedata
		.chrom_seg_23_s1_chipselect                    (mm_interconnect_0_chrom_seg_23_s1_chipselect),             //                                        .chipselect
		.chrom_seg_24_s1_address                       (mm_interconnect_0_chrom_seg_24_s1_address),                //                         chrom_seg_24_s1.address
		.chrom_seg_24_s1_write                         (mm_interconnect_0_chrom_seg_24_s1_write),                  //                                        .write
		.chrom_seg_24_s1_readdata                      (mm_interconnect_0_chrom_seg_24_s1_readdata),               //                                        .readdata
		.chrom_seg_24_s1_writedata                     (mm_interconnect_0_chrom_seg_24_s1_writedata),              //                                        .writedata
		.chrom_seg_24_s1_chipselect                    (mm_interconnect_0_chrom_seg_24_s1_chipselect),             //                                        .chipselect
		.chrom_seg_25_s1_address                       (mm_interconnect_0_chrom_seg_25_s1_address),                //                         chrom_seg_25_s1.address
		.chrom_seg_25_s1_write                         (mm_interconnect_0_chrom_seg_25_s1_write),                  //                                        .write
		.chrom_seg_25_s1_readdata                      (mm_interconnect_0_chrom_seg_25_s1_readdata),               //                                        .readdata
		.chrom_seg_25_s1_writedata                     (mm_interconnect_0_chrom_seg_25_s1_writedata),              //                                        .writedata
		.chrom_seg_25_s1_chipselect                    (mm_interconnect_0_chrom_seg_25_s1_chipselect),             //                                        .chipselect
		.chrom_seg_26_s1_address                       (mm_interconnect_0_chrom_seg_26_s1_address),                //                         chrom_seg_26_s1.address
		.chrom_seg_26_s1_write                         (mm_interconnect_0_chrom_seg_26_s1_write),                  //                                        .write
		.chrom_seg_26_s1_readdata                      (mm_interconnect_0_chrom_seg_26_s1_readdata),               //                                        .readdata
		.chrom_seg_26_s1_writedata                     (mm_interconnect_0_chrom_seg_26_s1_writedata),              //                                        .writedata
		.chrom_seg_26_s1_chipselect                    (mm_interconnect_0_chrom_seg_26_s1_chipselect),             //                                        .chipselect
		.chrom_seg_27_s1_address                       (mm_interconnect_0_chrom_seg_27_s1_address),                //                         chrom_seg_27_s1.address
		.chrom_seg_27_s1_write                         (mm_interconnect_0_chrom_seg_27_s1_write),                  //                                        .write
		.chrom_seg_27_s1_readdata                      (mm_interconnect_0_chrom_seg_27_s1_readdata),               //                                        .readdata
		.chrom_seg_27_s1_writedata                     (mm_interconnect_0_chrom_seg_27_s1_writedata),              //                                        .writedata
		.chrom_seg_27_s1_chipselect                    (mm_interconnect_0_chrom_seg_27_s1_chipselect),             //                                        .chipselect
		.chrom_seg_28_s1_address                       (mm_interconnect_0_chrom_seg_28_s1_address),                //                         chrom_seg_28_s1.address
		.chrom_seg_28_s1_write                         (mm_interconnect_0_chrom_seg_28_s1_write),                  //                                        .write
		.chrom_seg_28_s1_readdata                      (mm_interconnect_0_chrom_seg_28_s1_readdata),               //                                        .readdata
		.chrom_seg_28_s1_writedata                     (mm_interconnect_0_chrom_seg_28_s1_writedata),              //                                        .writedata
		.chrom_seg_28_s1_chipselect                    (mm_interconnect_0_chrom_seg_28_s1_chipselect),             //                                        .chipselect
		.chrom_seg_29_s1_address                       (mm_interconnect_0_chrom_seg_29_s1_address),                //                         chrom_seg_29_s1.address
		.chrom_seg_29_s1_write                         (mm_interconnect_0_chrom_seg_29_s1_write),                  //                                        .write
		.chrom_seg_29_s1_readdata                      (mm_interconnect_0_chrom_seg_29_s1_readdata),               //                                        .readdata
		.chrom_seg_29_s1_writedata                     (mm_interconnect_0_chrom_seg_29_s1_writedata),              //                                        .writedata
		.chrom_seg_29_s1_chipselect                    (mm_interconnect_0_chrom_seg_29_s1_chipselect),             //                                        .chipselect
		.chrom_seg_3_s1_address                        (mm_interconnect_0_chrom_seg_3_s1_address),                 //                          chrom_seg_3_s1.address
		.chrom_seg_3_s1_write                          (mm_interconnect_0_chrom_seg_3_s1_write),                   //                                        .write
		.chrom_seg_3_s1_readdata                       (mm_interconnect_0_chrom_seg_3_s1_readdata),                //                                        .readdata
		.chrom_seg_3_s1_writedata                      (mm_interconnect_0_chrom_seg_3_s1_writedata),               //                                        .writedata
		.chrom_seg_3_s1_chipselect                     (mm_interconnect_0_chrom_seg_3_s1_chipselect),              //                                        .chipselect
		.chrom_seg_30_s1_address                       (mm_interconnect_0_chrom_seg_30_s1_address),                //                         chrom_seg_30_s1.address
		.chrom_seg_30_s1_write                         (mm_interconnect_0_chrom_seg_30_s1_write),                  //                                        .write
		.chrom_seg_30_s1_readdata                      (mm_interconnect_0_chrom_seg_30_s1_readdata),               //                                        .readdata
		.chrom_seg_30_s1_writedata                     (mm_interconnect_0_chrom_seg_30_s1_writedata),              //                                        .writedata
		.chrom_seg_30_s1_chipselect                    (mm_interconnect_0_chrom_seg_30_s1_chipselect),             //                                        .chipselect
		.chrom_seg_4_s1_address                        (mm_interconnect_0_chrom_seg_4_s1_address),                 //                          chrom_seg_4_s1.address
		.chrom_seg_4_s1_write                          (mm_interconnect_0_chrom_seg_4_s1_write),                   //                                        .write
		.chrom_seg_4_s1_readdata                       (mm_interconnect_0_chrom_seg_4_s1_readdata),                //                                        .readdata
		.chrom_seg_4_s1_writedata                      (mm_interconnect_0_chrom_seg_4_s1_writedata),               //                                        .writedata
		.chrom_seg_4_s1_chipselect                     (mm_interconnect_0_chrom_seg_4_s1_chipselect),              //                                        .chipselect
		.chrom_seg_5_s1_address                        (mm_interconnect_0_chrom_seg_5_s1_address),                 //                          chrom_seg_5_s1.address
		.chrom_seg_5_s1_write                          (mm_interconnect_0_chrom_seg_5_s1_write),                   //                                        .write
		.chrom_seg_5_s1_readdata                       (mm_interconnect_0_chrom_seg_5_s1_readdata),                //                                        .readdata
		.chrom_seg_5_s1_writedata                      (mm_interconnect_0_chrom_seg_5_s1_writedata),               //                                        .writedata
		.chrom_seg_5_s1_chipselect                     (mm_interconnect_0_chrom_seg_5_s1_chipselect),              //                                        .chipselect
		.chrom_seg_6_s1_address                        (mm_interconnect_0_chrom_seg_6_s1_address),                 //                          chrom_seg_6_s1.address
		.chrom_seg_6_s1_write                          (mm_interconnect_0_chrom_seg_6_s1_write),                   //                                        .write
		.chrom_seg_6_s1_readdata                       (mm_interconnect_0_chrom_seg_6_s1_readdata),                //                                        .readdata
		.chrom_seg_6_s1_writedata                      (mm_interconnect_0_chrom_seg_6_s1_writedata),               //                                        .writedata
		.chrom_seg_6_s1_chipselect                     (mm_interconnect_0_chrom_seg_6_s1_chipselect),              //                                        .chipselect
		.chrom_seg_7_s1_address                        (mm_interconnect_0_chrom_seg_7_s1_address),                 //                          chrom_seg_7_s1.address
		.chrom_seg_7_s1_write                          (mm_interconnect_0_chrom_seg_7_s1_write),                   //                                        .write
		.chrom_seg_7_s1_readdata                       (mm_interconnect_0_chrom_seg_7_s1_readdata),                //                                        .readdata
		.chrom_seg_7_s1_writedata                      (mm_interconnect_0_chrom_seg_7_s1_writedata),               //                                        .writedata
		.chrom_seg_7_s1_chipselect                     (mm_interconnect_0_chrom_seg_7_s1_chipselect),              //                                        .chipselect
		.chrom_seg_8_s1_address                        (mm_interconnect_0_chrom_seg_8_s1_address),                 //                          chrom_seg_8_s1.address
		.chrom_seg_8_s1_write                          (mm_interconnect_0_chrom_seg_8_s1_write),                   //                                        .write
		.chrom_seg_8_s1_readdata                       (mm_interconnect_0_chrom_seg_8_s1_readdata),                //                                        .readdata
		.chrom_seg_8_s1_writedata                      (mm_interconnect_0_chrom_seg_8_s1_writedata),               //                                        .writedata
		.chrom_seg_8_s1_chipselect                     (mm_interconnect_0_chrom_seg_8_s1_chipselect),              //                                        .chipselect
		.chrom_seg_9_s1_address                        (mm_interconnect_0_chrom_seg_9_s1_address),                 //                          chrom_seg_9_s1.address
		.chrom_seg_9_s1_write                          (mm_interconnect_0_chrom_seg_9_s1_write),                   //                                        .write
		.chrom_seg_9_s1_readdata                       (mm_interconnect_0_chrom_seg_9_s1_readdata),                //                                        .readdata
		.chrom_seg_9_s1_writedata                      (mm_interconnect_0_chrom_seg_9_s1_writedata),               //                                        .writedata
		.chrom_seg_9_s1_chipselect                     (mm_interconnect_0_chrom_seg_9_s1_chipselect),              //                                        .chipselect
		.done_processing_chrom_s1_address              (mm_interconnect_0_done_processing_chrom_s1_address),       //                done_processing_chrom_s1.address
		.done_processing_chrom_s1_readdata             (mm_interconnect_0_done_processing_chrom_s1_readdata),      //                                        .readdata
		.done_processing_feedback_s1_address           (mm_interconnect_0_done_processing_feedback_s1_address),    //             done_processing_feedback_s1.address
		.done_processing_feedback_s1_write             (mm_interconnect_0_done_processing_feedback_s1_write),      //                                        .write
		.done_processing_feedback_s1_readdata          (mm_interconnect_0_done_processing_feedback_s1_readdata),   //                                        .readdata
		.done_processing_feedback_s1_writedata         (mm_interconnect_0_done_processing_feedback_s1_writedata),  //                                        .writedata
		.done_processing_feedback_s1_chipselect        (mm_interconnect_0_done_processing_feedback_s1_chipselect), //                                        .chipselect
		.error_sum_0_s1_address                        (mm_interconnect_0_error_sum_0_s1_address),                 //                          error_sum_0_s1.address
		.error_sum_0_s1_readdata                       (mm_interconnect_0_error_sum_0_s1_readdata),                //                                        .readdata
		.error_sum_1_s1_address                        (mm_interconnect_0_error_sum_1_s1_address),                 //                          error_sum_1_s1.address
		.error_sum_1_s1_readdata                       (mm_interconnect_0_error_sum_1_s1_readdata),                //                                        .readdata
		.error_sum_2_s1_address                        (mm_interconnect_0_error_sum_2_s1_address),                 //                          error_sum_2_s1.address
		.error_sum_2_s1_readdata                       (mm_interconnect_0_error_sum_2_s1_readdata),                //                                        .readdata
		.error_sum_3_s1_address                        (mm_interconnect_0_error_sum_3_s1_address),                 //                          error_sum_3_s1.address
		.error_sum_3_s1_readdata                       (mm_interconnect_0_error_sum_3_s1_readdata),                //                                        .readdata
		.error_sum_4_s1_address                        (mm_interconnect_0_error_sum_4_s1_address),                 //                          error_sum_4_s1.address
		.error_sum_4_s1_readdata                       (mm_interconnect_0_error_sum_4_s1_readdata),                //                                        .readdata
		.error_sum_5_s1_address                        (mm_interconnect_0_error_sum_5_s1_address),                 //                          error_sum_5_s1.address
		.error_sum_5_s1_readdata                       (mm_interconnect_0_error_sum_5_s1_readdata),                //                                        .readdata
		.error_sum_6_s1_address                        (mm_interconnect_0_error_sum_6_s1_address),                 //                          error_sum_6_s1.address
		.error_sum_6_s1_readdata                       (mm_interconnect_0_error_sum_6_s1_readdata),                //                                        .readdata
		.error_sum_7_s1_address                        (mm_interconnect_0_error_sum_7_s1_address),                 //                          error_sum_7_s1.address
		.error_sum_7_s1_readdata                       (mm_interconnect_0_error_sum_7_s1_readdata),                //                                        .readdata
		.expected_output_0_s1_address                  (mm_interconnect_0_expected_output_0_s1_address),           //                    expected_output_0_s1.address
		.expected_output_0_s1_write                    (mm_interconnect_0_expected_output_0_s1_write),             //                                        .write
		.expected_output_0_s1_readdata                 (mm_interconnect_0_expected_output_0_s1_readdata),          //                                        .readdata
		.expected_output_0_s1_writedata                (mm_interconnect_0_expected_output_0_s1_writedata),         //                                        .writedata
		.expected_output_0_s1_chipselect               (mm_interconnect_0_expected_output_0_s1_chipselect),        //                                        .chipselect
		.input_sequence_0_s1_address                   (mm_interconnect_0_input_sequence_0_s1_address),            //                     input_sequence_0_s1.address
		.input_sequence_0_s1_write                     (mm_interconnect_0_input_sequence_0_s1_write),              //                                        .write
		.input_sequence_0_s1_readdata                  (mm_interconnect_0_input_sequence_0_s1_readdata),           //                                        .readdata
		.input_sequence_0_s1_writedata                 (mm_interconnect_0_input_sequence_0_s1_writedata),          //                                        .writedata
		.input_sequence_0_s1_chipselect                (mm_interconnect_0_input_sequence_0_s1_chipselect),         //                                        .chipselect
		.nextSample_s1_address                         (mm_interconnect_0_nextsample_s1_address),                  //                           nextSample_s1.address
		.nextSample_s1_readdata                        (mm_interconnect_0_nextsample_s1_readdata),                 //                                        .readdata
		.preparingNextSample_s1_address                (mm_interconnect_0_preparingnextsample_s1_address),         //                  preparingNextSample_s1.address
		.preparingNextSample_s1_write                  (mm_interconnect_0_preparingnextsample_s1_write),           //                                        .write
		.preparingNextSample_s1_readdata               (mm_interconnect_0_preparingnextsample_s1_readdata),        //                                        .readdata
		.preparingNextSample_s1_writedata              (mm_interconnect_0_preparingnextsample_s1_writedata),       //                                        .writedata
		.preparingNextSample_s1_chipselect             (mm_interconnect_0_preparingnextsample_s1_chipselect),      //                                        .chipselect
		.ready_to_process_s1_address                   (mm_interconnect_0_ready_to_process_s1_address),            //                     ready_to_process_s1.address
		.ready_to_process_s1_readdata                  (mm_interconnect_0_ready_to_process_s1_readdata),           //                                        .readdata
		.sampleIndex_s1_address                        (mm_interconnect_0_sampleindex_s1_address),                 //                          sampleIndex_s1.address
		.sampleIndex_s1_write                          (mm_interconnect_0_sampleindex_s1_write),                   //                                        .write
		.sampleIndex_s1_readdata                       (mm_interconnect_0_sampleindex_s1_readdata),                //                                        .readdata
		.sampleIndex_s1_writedata                      (mm_interconnect_0_sampleindex_s1_writedata),               //                                        .writedata
		.sampleIndex_s1_chipselect                     (mm_interconnect_0_sampleindex_s1_chipselect),              //                                        .chipselect
		.sequences_to_process_s1_address               (mm_interconnect_0_sequences_to_process_s1_address),        //                 sequences_to_process_s1.address
		.sequences_to_process_s1_write                 (mm_interconnect_0_sequences_to_process_s1_write),          //                                        .write
		.sequences_to_process_s1_readdata              (mm_interconnect_0_sequences_to_process_s1_readdata),       //                                        .readdata
		.sequences_to_process_s1_writedata             (mm_interconnect_0_sequences_to_process_s1_writedata),      //                                        .writedata
		.sequences_to_process_s1_chipselect            (mm_interconnect_0_sequences_to_process_s1_chipselect),     //                                        .chipselect
		.start_processing_chrom_s1_address             (mm_interconnect_0_start_processing_chrom_s1_address),      //               start_processing_chrom_s1.address
		.start_processing_chrom_s1_write               (mm_interconnect_0_start_processing_chrom_s1_write),        //                                        .write
		.start_processing_chrom_s1_readdata            (mm_interconnect_0_start_processing_chrom_s1_readdata),     //                                        .readdata
		.start_processing_chrom_s1_writedata           (mm_interconnect_0_start_processing_chrom_s1_writedata),    //                                        .writedata
		.start_processing_chrom_s1_chipselect          (mm_interconnect_0_start_processing_chrom_s1_chipselect),   //                                        .chipselect
		.two_port_mem_s1_address                       (mm_interconnect_0_two_port_mem_s1_address),                //                         two_port_mem_s1.address
		.two_port_mem_s1_write                         (mm_interconnect_0_two_port_mem_s1_write),                  //                                        .write
		.two_port_mem_s1_readdata                      (mm_interconnect_0_two_port_mem_s1_readdata),               //                                        .readdata
		.two_port_mem_s1_writedata                     (mm_interconnect_0_two_port_mem_s1_writedata),              //                                        .writedata
		.two_port_mem_s1_byteenable                    (mm_interconnect_0_two_port_mem_s1_byteenable),             //                                        .byteenable
		.two_port_mem_s1_chipselect                    (mm_interconnect_0_two_port_mem_s1_chipselect),             //                                        .chipselect
		.two_port_mem_s1_clken                         (mm_interconnect_0_two_port_mem_s1_clken),                  //                                        .clken
		.two_port_mem_correct_s1_address               (mm_interconnect_0_two_port_mem_correct_s1_address),        //                 two_port_mem_correct_s1.address
		.two_port_mem_correct_s1_write                 (mm_interconnect_0_two_port_mem_correct_s1_write),          //                                        .write
		.two_port_mem_correct_s1_readdata              (mm_interconnect_0_two_port_mem_correct_s1_readdata),       //                                        .readdata
		.two_port_mem_correct_s1_writedata             (mm_interconnect_0_two_port_mem_correct_s1_writedata),      //                                        .writedata
		.two_port_mem_correct_s1_byteenable            (mm_interconnect_0_two_port_mem_correct_s1_byteenable),     //                                        .byteenable
		.two_port_mem_correct_s1_chipselect            (mm_interconnect_0_two_port_mem_correct_s1_chipselect),     //                                        .chipselect
		.two_port_mem_correct_s1_clken                 (mm_interconnect_0_two_port_mem_correct_s1_clken),          //                                        .clken
		.valid_output_0_s1_address                     (mm_interconnect_0_valid_output_0_s1_address),              //                       valid_output_0_s1.address
		.valid_output_0_s1_write                       (mm_interconnect_0_valid_output_0_s1_write),                //                                        .write
		.valid_output_0_s1_readdata                    (mm_interconnect_0_valid_output_0_s1_readdata),             //                                        .readdata
		.valid_output_0_s1_writedata                   (mm_interconnect_0_valid_output_0_s1_writedata),            //                                        .writedata
		.valid_output_0_s1_chipselect                  (mm_interconnect_0_valid_output_0_s1_chipselect),           //                                        .chipselect
		.writeSample_s1_address                        (mm_interconnect_0_writesample_s1_address),                 //                          writeSample_s1.address
		.writeSample_s1_write                          (mm_interconnect_0_writesample_s1_write),                   //                                        .write
		.writeSample_s1_readdata                       (mm_interconnect_0_writesample_s1_readdata),                //                                        .readdata
		.writeSample_s1_writedata                      (mm_interconnect_0_writesample_s1_writedata),               //                                        .writedata
		.writeSample_s1_chipselect                     (mm_interconnect_0_writesample_s1_chipselect)               //                                        .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
